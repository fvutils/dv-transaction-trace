
package dvtt;
    int _dvtt_debug_level = 0;

endpackage

